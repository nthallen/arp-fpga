--
-- VHDL Architecture idx_fpga_lib.ana_ram.beh
--
-- Created:
--          by - nort.UNKNOWN (NORT-NBX200T)
--          at - 10:00:43 10/14/2010
--
-- using Mentor Graphics HDL Designer(TM) 2009.2 (Build 10)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
Library UNISIM;
use UNISIM.vcomponents.all;

ENTITY ana_ram IS
  PORT (
    RD_ADDR : IN std_logic_vector(7 DOWNTO 0);
    WR_ADDR : IN std_logic_vector(7 DOWNTO 0);
    RD_DATA : OUT std_logic_vector(31 DOWNTO 0);
    WR_DATA : IN std_logic_vector(31 DOWNTO 0);
    WREN : IN std_ulogic;
    RDEN : IN std_ulogic;
    CLK : IN std_ulogic;
    RST : IN std_ulogic
  );
END ENTITY ana_ram;

--
ARCHITECTURE beh OF ana_ram IS
  SIGNAL DOPADOP : std_logic_vector(1 downto 0);
  SIGNAL DOPBDOP : std_logic_vector(1 downto 0);
  SIGNAL ADDRAWRADDR : std_logic_vector(12 downto 0);
  SIGNAL ADDRBRDADDR : std_logic_vector(12 downto 0);
  SIGNAL DIPADIP : std_logic_vector(1 downto 0);
  SIGNAL DIPBDIP : std_logic_vector(1 downto 0);
  SIGNAL WEAWEL : std_logic_vector(1 downto 0);
  SIGNAL WEBWEU : std_logic_vector(1 downto 0);

  COMPONENT RAMB8BWER is
    generic (
      DATA_WIDTH_A : integer := 0;
      DATA_WIDTH_B : integer := 0;
      DOA_REG : integer := 0;
      DOB_REG : integer := 0;
      EN_RSTRAM_A : boolean := TRUE;
      EN_RSTRAM_B : boolean := TRUE;
      INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_A : bit_vector := X"00000";
      INIT_B : bit_vector := X"00000";
      INIT_FILE : string := "NONE";
      RAM_MODE : string := "TDP";
      RSTTYPE  : string := "SYNC";
      RST_PRIORITY_A : string := "SR";
      RST_PRIORITY_B : string := "SR";
      SETUP_ALL : time := 1000 ps;
      SETUP_READ_FIRST : time := 3000 ps;
      SIM_COLLISION_CHECK : string := "ALL";
      SRVAL_A : bit_vector := X"00000";
      SRVAL_B : bit_vector := X"00000";
      WRITE_MODE_A : string := "WRITE_FIRST";
      WRITE_MODE_B : string := "WRITE_FIRST"
      );

    port (

      DOADO : out std_logic_vector(15 downto 0);
      DOBDO : out std_logic_vector(15 downto 0);
      DOPADOP : out std_logic_vector(1 downto 0);
      DOPBDOP : out std_logic_vector(1 downto 0);

      ADDRAWRADDR : in std_logic_vector(12 downto 0);
      ADDRBRDADDR : in std_logic_vector(12 downto 0);
      CLKAWRCLK : in std_ulogic;
      CLKBRDCLK : in std_ulogic;
      DIADI : in std_logic_vector(15 downto 0);
      DIBDI : in std_logic_vector(15 downto 0);
      DIPADIP : in std_logic_vector(1 downto 0);
      DIPBDIP : in std_logic_vector(1 downto 0);
      ENAWREN : in std_ulogic;
      ENBRDEN : in std_ulogic;
      REGCEA : in std_ulogic;
      REGCEBREGCE : in std_ulogic;
      RSTA : in std_ulogic;
      RSTBRST : in std_ulogic;
      WEAWEL : in std_logic_vector(1 downto 0);
      WEBWEU : in std_logic_vector(1 downto 0)

      ); 
  end component;

BEGIN

   -- RAMB8BWER: 8K-bit Data and 1K-bit Parity Configurable Synchronous Block RAM
   --            Spartan-6
   -- Xilinx HDL Language Template, version 12.1

   RAMB8BWER_inst : RAMB8BWER
   generic map (
      -- DATA_WIDTH_A/DATA_WIDTH_B: If RAM_MODE=TDP: 0, 1, 2, 4, 9 or 18; If RAM_MODE=SDP: 36
      DATA_WIDTH_A => 36,
      DATA_WIDTH_B => 36,
      -- DOA_REG/DOB_REG: Optional output register (0 or 1)
      DOA_REG => 0,
      DOB_REG => 0,
      -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
      EN_RSTRAM_A => TRUE,
      EN_RSTRAM_B => TRUE,
      -- INITP_00 to INITP_03: Initial memory contents.
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- INIT_00 to INIT_1F: Initial memory contents.
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- INIT_A/INIT_B: Initial values on output port
      INIT_A => X"00000",
      INIT_B => X"00000",
      -- INIT_FILE: Optional file used to specify initial RAM contents
      INIT_FILE => "NONE",
      -- RAM_MODE: "SDP" or "TDP" 
      RAM_MODE => "SDP",
      -- RSTTYPE: "SYNC" or "ASYNC" 
      RSTTYPE => "SYNC",
      -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
      RST_PRIORITY_A => "CE",
      RST_PRIORITY_B => "CE",
      -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
      SIM_COLLISION_CHECK => "ALL",
      -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
      SRVAL_A => X"00000",
      SRVAL_B => X"00000",
      -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
      WRITE_MODE_A => "READ_FIRST",
      WRITE_MODE_B => "READ_FIRST" 
   )
   port map (
      DOADO => RD_DATA(15 DOWNTO 0),             -- 16-bit A port data/LSB data output
      DOBDO => RD_DATA(31 DOWNTO 16),             -- 16-bit B port data/MSB data output
      DOPADOP => DOPADOP,         -- 2-bit A port parity/LSB parity output
      DOPBDOP => DOPBDOP,         -- 2-bit B port parity/MSB parity output
      ADDRAWRADDR => ADDRAWRADDR, -- 13-bit A port address/Write address input
      ADDRBRDADDR => ADDRBRDADDR, -- 13-bit B port address/Read address input
      CLKAWRCLK => CLK,           -- 1-bit A port clock/Write clock input
      CLKBRDCLK => CLK,           -- 1-bit B port clock/Read clock input
      DIADI => WR_DATA(15 DOWNTO 0),  -- 16-bit A port data/LSB data input
      DIBDI => WR_DATA(31 DOWNTO 16), -- 16-bit B port data/MSB data input
      DIPADIP => DIPADIP,         -- 2-bit A port parity/LSB parity input
      DIPBDIP => DIPBDIP,         -- 2-bit B port parity/MSB parity input
      ENAWREN => WREN,            -- 1-bit A port enable/Write enable input
      ENBRDEN => RDEN,            -- 1-bit B port enable/Read enable input
      REGCEA => '0',              -- 1-bit A port register enable input
      REGCEBREGCE => '0',         -- 1-bit B port register enable/Register enable input
      RSTA => RST,                -- 1-bit A port set/reset input
      RSTBRST => RST,             -- 1-bit B port set/reset input
      WEAWEL => WEAWEL,           -- 2-bit A port write enable input
      WEBWEU => WEBWEU            -- 2-bit B port write enable input
   );

  ADDRAWRADDR(12 DOWNTO 5) <= WR_ADDR;
  ADDRAWRADDR(4 DOWNTO 0) <= (others => '0');
  ADDRBRDADDR(12 DOWNTO 5) <= RD_ADDR;
  ADDRBRDADDR(4 DOWNTO 0) <= (others => '0');
  DIPADIP <= (others => '0');
  DIPBDIP <= (others => '0');
  WEAWEL(1) <= WREN;
  WEAWEL(0) <= WREN;
  WEBWEU(1) <= WREN;
  WEBWEU(0) <= WREN;
END ARCHITECTURE beh;

