--
-- VHDL Architecture idx_fpga_lib.ana_ram.beh
--
-- Created:
--          by - nort.UNKNOWN (NORT-NBX200T)
--          at - 10:00:43 10/14/2010
--
-- using Mentor Graphics HDL Designer(TM) 2009.2 (Build 10)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
Library unimacro;
USE unimacro.VCOMPONENTS.all;

ENTITY ana_ram IS
  PORT (
    RD_ADDR : IN std_logic_vector(7 DOWNTO 0);
    WR_ADDR : IN std_logic_vector(7 DOWNTO 0);
    RD_DATA : OUT std_logic_vector(31 DOWNTO 0);
    WR_DATA : IN std_logic_vector(31 DOWNTO 0);
    WREN : IN std_ulogic_vector(1 DOWNTO 0);
    RDEN : IN std_ulogic;
    OE : IN std_ulogic;
    CLK : IN std_ulogic;
    RST : IN std_ulogic
  );
END ENTITY ana_ram;

ARCHITECTURE beh OF ana_ram IS
  SIGNAL WREN_int : std_ulogic;
  SIGNAL RDEN_int : std_ulogic;
  SIGNAL WE : std_logic_vector(3 DOWNTO 0);
  SIGNAL RD_DATA_int : std_logic_vector(31 DOWNTO 0);
  SIGNAL RDEN_dly : std_ulogic;
  SIGNAL RAM_RD_ADDR : std_logic_vector(8 DOWNTO 0);
  SIGNAL RAM_WR_ADDR : std_logic_vector(8 DOWNTO 0);

  COMPONENT BRAM_SDP_MACRO is
  generic (
      BRAM_SIZE : string := "18Kb";
      DEVICE : string := "VIRTEX5";
      DO_REG : integer := 0;
      INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_40 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_41 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_42 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_43 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_44 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_45 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_46 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_47 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_48 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_49 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_4A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_4B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_4C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_4D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_4E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_4F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_50 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_51 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_52 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_53 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_54 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_55 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_56 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_57 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_58 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_59 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_5A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_5B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_5C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_5D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_5E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_5F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_60 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_61 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_62 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_63 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_64 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_65 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_66 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_67 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_68 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_69 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_6A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_6B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_6C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_6D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_6E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_6F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_70 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_71 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_72 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_73 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_74 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_75 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_76 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_77 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_78 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_79 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_7A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_7B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_7C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_7D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_7E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_7F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT : bit_vector := X"000000000000000000";
      INIT_FILE : string := "NONE";
      READ_WIDTH : integer := 0;
      WRITE_WIDTH : integer := 0;
      SIM_COLLISION_CHECK : string := "ALL";
      SIM_MODE : string := "SAFE"; -- This parameter is valid only for Virtex5
      SRVAL : bit_vector := X"000000000000000000"
    );
  -- ports are unconstrained arrays
  port (
    
      DO : out std_logic_vector;

      DI : in std_logic_vector;
      RDADDR : in std_logic_vector;
      RDCLK : in std_ulogic;
      RDEN : in std_ulogic;
      REGCE : in std_ulogic;
      RST : in std_ulogic;
      WE : in std_logic_vector;
      WRADDR : in std_logic_vector;
      WRCLK : in std_ulogic;
      WREN : in std_ulogic

    );
  end COMPONENT;

  FOR ALL : bram_sdp_macro USE ENTITY unimacro.bram_sdp_macro;
BEGIN
  bram_sdp_macro_inst : bram_sdp_macro
  generic map (
     BRAM_SIZE => "18Kb", -- Target BRAM, "18Kb" or "36Kb"
     DEVICE => "SPARTAN6", -- Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
     WRITE_WIDTH => 32,    -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
     READ_WIDTH => 32,     -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
     DO_REG => 0, -- Optional output register (0 or 1)
     INIT_FILE => "NONE",
     SIM_COLLISION_CHECK => "ALL", -- Collision check enable "ALL", "WARNING_ONLY", 
                                   -- "GENERATE_X_ONLY" or "NONE"       
     SIM_MODE => "SAFE", -- Simulation: "SAFE" vs "FAST", 
                         -- see "Synthesis and Simulation Design Guide" for details
     SRVAL => X"000000000000000000", --  Set/Reset value for port output
     INIT => X"000000000000000000", --  Initial values on output port
     -- The following INIT_xx declarations specify the initial contents of the RAM
     INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
     
     -- The next set of INIT_xx are valid when configured as 36Kb
     INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
     INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
     
     -- The next set of INITP_xx are for the parity bits
     INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
     
     -- The next set of INIT_xx are valid when configured as 36Kb
     INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
     INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
     DO => RD_DATA_int, -- Output read data port
     DI => WR_DATA,     -- Input write data port
     RDADDR => RAM_RD_ADDR, -- Input read address
     RDCLK => CLK,      -- Input read clock
     RDEN => RDEN_int,  -- Input read port enable
     REGCE => '0',    -- Input read output register enable
     RST => RST,        -- Input reset 
     WE => WE,          -- Input write enable
     WRADDR => RAM_WR_ADDR, -- Input write address
     WRCLK => CLK,      -- Input write clock
     WREN => WREN_int   -- Input write port enable
  );
  
  RAM_RD_ADDR <= '0' & RD_ADDR;
  RAM_WR_ADDR <= '0' & WR_ADDR;

  Wr_En : Process (WREN) IS
  Begin
    if WREN = "11" then
      WREN_int <= '1';
    else
      WREN_int <= '0';
    end if;
  End Process;

  Rd_En : Process ( CLK, RST, RDEN, RDEN_dly ) IS
  Begin
    if RST = '1' then
      RDEN_dly <= '0';
    elsif CLK'Event AND CLK = '1' then
      RDEN_dly <= RDEN;
    end if;
    if RDEN = '1' AND RDEN_dly = '0' then
      RDEN_int <= '1';
    else
      RDEN_int <= '0';
    end if;
  End Process;
  
  Out_En : Process (OE,RD_DATA_int) Is
  Begin
    if OE = '1' then
      RD_DATA <= RD_DATA_int;
    else
      RD_DATA <= (others => 'Z');
    end if;
  End Process;

  WE(0) <= WREN_int;
  WE(1) <= WREN_int;
  WE(2) <= WREN_int;
  WE(3) <= WREN_int;
End Architecture beh;

